%@ Swedish hyphenation patterns.
%
% Copyright (c) 2014 - 2018 Steffen (Daode) Nurpmeso <steffen@sdaoden.eu>.
%
% Copyright 1994 by Jan Michael Rynning. All rights reserved.
%
% This program may be distributed and/or modified under the conditions of
% the LaTeX Project Public License, either version 1.2 of this license or
% (at your option) any later version.  The latest version of this license
% is in http://www.latex-project.org/lppl.txt and version 1.2 or later is
% part of all distributions of LaTeX version 1999/12/01 or later.
%
% Last update: 1994-03-03 (March 3, 1994).
% Revision history:
% 1991-01-08: First version available for anonymous FTP.
% 1991-08-08: Changed \aa to \aa0 at end of line, to stop TeX from
%             concatenating the patterns.
% 1991-09-03: Cleaned up lots of inconsistencies in the dictionary.
%             As a consequence, the patterns shrunk a lot.  Also
%             added some 4000 one-syllable words, some of which were
%             hyphenated by the old patterns, and some 1500 compound
%             words, about half of which were incorrectly hyphenated
%             by the old patterns.
% 1991-11-01: Added another some 6200 compound words, all of which were
%             incorrectly hyphenated by the old patterns.
% 1991-11-13: Added another some 6500 compound words, all of which were
%             incorrectly hyphenated by the old patterns.
% 1992-01-30: Changed macros to ^^, for use with LaTeX and dc fonts.
% 1994-03-03: The hyphenated dictionary now contains about 118,000 words.
%             The hyphenation now works much better for compound words.
%             Patgen parameters: 1 2 20, 2 1 8, 1 4 7, 3 2 1, 1 10000 4.
%
% This file contains Swedish hyphenation patterns for TeX.  It assumes
% that you have fonts with the Swedish letters in the positions where
% they occur in ISO Latin 1 (ISO 8859/1):
% Letter:   \AA  \"A  \"O  \'E  \aa  \"a  \"o  \'e
% Position: "C5  "C4  "D6  "C9  "E5  "E4  "F6  "E9
%
% Load this file into initex after plain.tex (or lplain.tex, splain.tex,
% or whatever).
%
% The patterns were generated in such a way that they will hyphenate
% correctly if \lefthyphenmin>=1 and \righthyphenmin>=2.
%
% These hyphenation patterns work quite well for simple words, but not
% quite as well for compound words.  I'm working on improving the quality,
% by adding more words.  If you know any Swedish words which are not
% correctly hypheneted using these patterns, or if you have questions or
% comments, please contact me:
%
% Jan Michael Rynning <jmr@incolumitas.se>
% --------------------------------------------------------------------------
\message{Swedish hyphenation patterns, Jan Michael Rynning, 1994-03-03.}
{
% Set \catcode, \uccode, and \lccode for the Swedish letters.
% This should be done for all letters, really.
\catcode`^^c5=11 \catcode`^^c4=11 \catcode`^^d6=11 \catcode`^^c9=11
\catcode`^^e5=11 \catcode`^^e4=11 \catcode`^^f6=11 \catcode`^^e9=11
\uccode`^^c5=`^^c5 \uccode`^^c4=`^^c4 \uccode`^^d6=`^^d6 \uccode`^^c9=`^^c9
\uccode`^^e5=`^^c5 \uccode`^^e4=`^^c4 \uccode`^^f6=`^^d6 \uccode`^^e9=`^^c9
\lccode`^^c5=`^^e5 \lccode`^^c4=`^^e4 \lccode`^^d6=`^^f6 \lccode`^^c9=`^^e9
\lccode`^^e5=`^^e5 \lccode`^^e4=`^^e4 \lccode`^^f6=`^^f6 \lccode`^^e9=`^^e9
\patterns{ % just type <return> if you're not using INITEX
.a4b
.ab5i
.ab5ol
.ab3r
.ac3
.a4d
.a3dr
.ad3s
.a5g4ra
.a5gre
.a5kl
.a5le
.al4pr
.a3lu
.am4br
.amp3l
.a5mu
.and4rar
.a2n5es
.ang4er
.an5go
.an5s
.ap1p
.as2k
.a3sket
.as4t
.a5sten
.a3sti
.a5ta
.at3t
.au3st
.a4val
.av3s4
.b4
.bak5s
.ben5s
.bild3s
.bo2k
.bort1
.cis4
.cy5klop
.d4
.d^^e4r3
.ek1v
.e3l4a
.e2l5in
.en5st
.e4n^^e4
.e2r3i
.e2s
.e5skad
.es3kal
.es5kap
.es4t
.e5strad
.e3tr
.evan5
.ex3
.f4
.feb3r
.fram3
.fres5
.f^^e5gel3
.f^^f6r1a
.f^^f6r1en
.g2
.gu4l^^e4
.gus3
.he2m
.hu5sa
.ib4
.ik4
.im3p
.i2n1
.i4na
.in3d
.in4ger
.ink2
.in3s2
.in3t
.is5ka
.i3so
.k4
.kans4k
.ko5li
.kort5s
.kring3
.krings2
.k^^f6p5s
.l2
.lak5r
.lek5tr
.lu2st
.m2
.mas2ke
.ma5skeri
.me4re
.minis4
.mj^^f6lk5s
.mon2s
.m^^e5n3s
.m^^e54st
.m^^e4n5sko
.m^^f6rk5r
.n4
.ner1
.no4n
.n^^f6d5r
.oc1ku
.ok3t
.o3kv
.o2ma
.o2mo
.om3s4
.o3mu
.on4k
.o3o
.ord3s
.o5sc
.o1s4k
.o3sl
.o3stra
.o3sv
.o3tr
.o1u
.p4
.papp5s
.pa3ste
.pa5sti
.pi5sti
.pres2s
.pub3lika
.r2
.re4gr
.re2ste
.runs4
.rym2d
.r^^f6ve5
.s4
.sa2k
.seg3r
.si5o
.sj^^f61
.sk4
.skott3s
.slut3s
.st4
.sta2m
.sten3s
.string4
.sup3p
.t4
.ta3bl
.ta4k
.tak5l
.tes3ta
.tig3r
.til4l
.ti3o
.topp5s
.tred2s
.tre3s
.tr^^e45k
.u3k
.ult5r
.ung2e
.up2
.u4ra
.ur3s
.u2t1
.u4ta
.u5trer
.ut5s
.v2
.var4t
.vatten3
.ved5s
.v^^e42g
.v^^e4g3s
.x2
.y2a
.y4e
.^^e5ng3
.^^e5r4s5
.^^e53st
.^^e5ter1
.^^e43ro
.^^f63ro
a2b
ab4bu
a5be
abel4s
abe2s
ab1l
ab3la
ab3ort
ab5ric
ab3rio
ab4sc
ab4sk
a5bu
ac4kes
ac4kis
ack3sk
ack3u4p
a5dag
a5dek
a5del
ad5ep
ad3j
ad3op
a5dran
a3dre
1adres
ad3ril
ad3ru
ad2s
a5ed
af4fo
3aff^^e4
1af3ri
af4tor
a1ga
aga4ra
a1ge
a2ge.
ag1gr
ag1l
ag5ord
ag3ro
a4gur
a4hj
aib4
a3iv
a1j
a3ka
a4kart
a5ke
a1ki
ak3n
a1ko
ak5ram
akri5s
ak3rob
ak4sta
1aktig
ak3tri
a1ku
a5kvari
ak3ve
a5k^^e5r
ak5^^e5t
4ak^^f6
a1la
al5adm
ali2br
a2lin
a5lin.
a3line
al3ins
ali5stik
a4lj
alk3ak
al2kv
al4k^^e4
all3st
al3l^^e5
alms4k
a1lo
al5ort
als5pa
al3tr
al4tu
al4t^^e4
a1lu
alu5s
alv3s
a1ly
a4maf
am4i
am4pr
am1s
am3^^e5t
a3m^^f6
ana4bo
an3alf
an3ark
an3c
anci5
an5dak
andel2s
an4dun
an4d^^e4n
a4nef
ang4es
an3gi
an1gr
aniu4
ank3r
ano2i
a4nok
a4nop
an5sce
ansis3t
an4sj
ans5ku
ans3li
ans3par
an1st
an4sto
an4sty
1ansvar
an4tj
an4tre
a1nu
a5ny
a3n^^f6
a1o
a1pe
a2pe.
ape4n3
a1pi
ap4lan
apo3str
1appara
apps4k
ap3ric
ap3rif
a5pris
ap2s
ap3se
aps5l
aps3p
apu5s
a5py
a5p^^e4
2ara
a4rann
a4rarv
1arb
4arbi
2arbo
4arbr
ar3dr
ard5st
a4rend
arg5si
2arh
a1ri
a4rigen
ar3ka
ark3lan
ar5kr
4arl
4arn.
ar4nal
a1ro
a2rob
4arp
ar2sa
ar5skal
arsk5l
ar2sv
ar4tro
arts5p
ar4tur
4aru
a4rur
a5rus
ar4v^^e4g
a3ry
a3r^^e4
2asa
asbe4
a1sc
as2h
asis5t
as3kis
a2sko
a4skr
as3ku
as5l
as3pa
as3pig
as2sk
as2s5op
as2sp
as2st
ass5up
as3ta
a5stard
as5ter
as5tiker
asti5o
as3to
as4tr
ast5rak
a5stral
ast3rol
as5t^^f6r
a3su
a4sul
a4sund
as2ut
as3v
a1sy
a2s5^^e5
a2s^^f6
a1t
ata5ra
a5te
ati5^^f6
a4tj
a2tr
a3tral
4atrar
a4t3re
at3ria
a3tric
at3rie
a5trik
a3tris
a3t4ro
a4tro.
at4ska
1attac
at2tak
at4tj
at4tos
att3s
a4tung
2au
au5b
au2t5a
3autom
aut5s
2a1va
a4vart
1avg
2a1vi
av3r
4a3v^^e4
a5^^e5
1b2
3ba
ba4di
ba4do
bad3s4
bak5l
ba4ko
ba4ku
bank5l
bas4ta
ba5stu
4bb
b4bak
b4batt
bbb4
bb3l
bb4ler
b4b3r
bb4so
4b3d
3be
be3d4r
be5e
be1k
4beld
be5lu
be3ly
be3l^^e5
be5l^^f6
beng4
be3n^^e5
be1r^^f6
be1s
be3sl
bes5s
be4sta
be4ste
be5su
be3tr
be3tv
be3u
4bex
2b3f
2b5h
3bi
bi3d4
4binv
bis3ko
bi5skv
b3je
b3k
b5lar
b5lat
ble4mo
b5len
5blera
3bles
5blid
3blikr
3bliks
4b3m
2b3n
3bo
bo4gr
bo2kl
bo1mu
5bon
bors5te
bor4ti
bort3r
borts2
bort3sl
bo1s
bo4sc
boy5
4b3p
2b5raf
4brar
2b5rati
3brik.
b3rika
3brike
3briks
b5rik^^f6
bru4st
3bry
3br^^f6
4b3s
b5sce
bs3ch
b4slan
b4sof
b4sp
bst4
b4stj
4b3t
3bu
bund4s
bus2st
b3v
3by
by5r
3b^^e5
b^^e5ng3
b^^e5t2s
3b^^e4
3b^^f6
b^^f6r2s
c2
5cap
c3c
1c4e
cens3t
3centr
ceu4s
4ch.
3chau
3chef
5choc
4cht
ch^^e4s3
ch^^f6r4
1ci
ci4lu
cim2
cipp4
4ck
c3ka
c3ke
c3ki
ck5j
ck1l
ck5lis
ck3n
c3ko
c4kordn
ck3org
c4kort
ck3r
ck4re
ck3sla
ckus2
ck3va
ck3ve
ck3v^^e4
ck5^^e4
ck3^^f6
cle2a
co2a
co4m
4cr
cros2
4cs
1cy
1d
3da
5da.
4dadr
dags3
2dak
5dako
da3li
5dam
da3m^^e5
4dand.
4d1ap
4darb
4dart
da4tr
dat5t
4dax
2db
4dc
dcen3
2dd
ddd4
ddi4s
d3dj
d4dos
dd3ra
dd3re
dd3ri
d3dr^^e4
dd2s
dds3v
3d2e
de1k4
4deko
4deld
del2sa
dels5ti
de5lut
d4en
denti5^^f6
den2to
de3pr
5der
der1k
de2ro
de5rol
der5sti
de4ru
de2s
de3se
de3sp
des3ti
d4et
de3tr
4dex
2d1f
df^^f63ra
2d1g
d3gl
2d5h
3di
dias4
di5el
di2gr
di3ka
di5ku
4dinf
din3g4o
4dinr
4dins
2dinsp
4dint
di1o
di4od
di3sc
di4sj
dis3ko
dis1kr
dis1p
dis5to
dis3tra
di4tre
2dj
d3jor
djup5p
3djur
2d3k2
4d5l
2d1m
2d1n
3do
d2ol
do5lo
4domr
dom2sk
5don
do4pak
4d5ord
4dori
4dort
d5ost
do3y
2d1p
2d2r2
d3rad
3d4rag
d3rand
d5rarb
d5rassera
d5ratu
3drej
d3ren
5dres
d3ret
d4ric
3drif
d3rig
4d5rik
d3rin
3d4riv
d5roc
3dropp
d3ror
4drot
drotts3
d3r^^e4kn
3dr^^e4kt
5dr^^e4n
d3r^^e4t
d5r^^f6d
4ds
d2s1an
d2se
ds5enh
d4sf
d2si
ds3ins
d2sj
dsk2
d3skef
ds4ken
d3ski
ds3kl
ds5kn
ds1l
ds4lot
ds4mo
d4sm^^e5
ds5n^^e5
d2so
ds3pl
ds3s4
ds3tal
d5stat
ds4te
dste4a
d5stig
ds3tin
ds5tro
d2su
ds1v
d2s^^f6
2d3t
3du
dub3ble
4dup
du1s
du2sc
du4ste
du5s^^f6
4dut
du4vu
2d1v
d3vr
2d3w
3dy
dy4kan
dy4ro
4dz
5d^^e5g
2d^^e5s
4d^^e5t
4d^^e4g
d^^e42r
3d^^f6
d^^f6ds1
4d^^f6g
4d^^f6p
d5^^f6st
d^^e94
e1a
e2ake
e4am
4eb
e2br
eb3ril
4ec
e3ch
echiff5
ecis4
e3co
e2d
e4dans
edd4r
edi4u
ed3j
e5dral
ed1sk
ed2sko
ed3s2l
edso4
e3d^^e5
e1e
e2ed
e4ei
ee2k5
e4en.
e4ene
e1f
ef4s
3efte
e1g
e3ga
e3ge
ege2l
eg1l
eg2ler
e3glera
e5gleri
e4gran
eg5rat
eg3rin
e5gru
egs3
e5g^^e5
eig2
ei5gn
e3ik
e1in
ei5sh
e1isk
e1jo
e3ju
e3j^^e4
e5j^^f6
e3ka
e1ki
e1kl
ek3lat
ek4le
ek3n
e1ko
ekord5s
ek3orr
ek4ret.
ek5ro
e1ku
e1kve
ek5vis
e1ky
e1k^^e4
e1la
el1akt
el4arb
3eld.
eleb3r
elekt3ri
el4fra
eli5ku
el3k4
el3li
ell3s
el3l^^e4
e1lo
e4lob
el3p
el2si
el5ug
e5luv
2e1l^^e4
e1m
e5mat
e5mis
emon1s
em5ort
emp5le
en5art
e2nav
en4ce
e4ned
e4nek
ene3r^^f6
2enj
en5klo
en3kn
en5kr
en5k^^e4
enning5
ennings2
eno2m
en3si
ens5ke
ens2m
en2sp
ens4te
ens4vin
en4s^^e5
ent4ha
en2t1r
ent4rat.
ent3rati
ent3ri
ent5ru
e5nus
2eny
2e1n^^e4
e1o
e2og
eo4i
e5or
2ep
e1pe
e1pi
e3pla
ep5le
epp2s3
epps5t
e1pr
ep3s
ep4tr
epu3b
e3p^^e5
er1ak
4eras
er3d4
erg4l
er4gu
er4g^^e5s
e1ri
e5rib
e4rinf
erings3
eri5stik
erk4lin
erl^^e44
er5na
e1ro
e3rob
e2rom
erp4
er3ra
er5sc
ers4ken
er3sl
ers4le
er4sta
er2ste
er3str
er3sv
e1ru
e5rum
e3ry
e5r^^e5d
e1r^^e4
e2sal
es5all
es3arm
e1sc
2ese
es4hi
esi4u
es2k
e4skan
es5kar
e4s3ken
es3ker
es5kul
e1sl
e5slag
es2mi
e1sp
es3pl
es2sk
ess5l^^e4
es2st
e3stal
es5ten.
esti2ge
es3tin
es5tor.
es4tr
est5rer
e3stru
est4r^^f6
e3st^^e5
es2u
e1sy
eta3b
e5ti
eti3^^f6
e1to
e5tri.
et3ris
e5tr^^e4
et2s
ets2ad
ets3kr
ets1l
ets3m
ets5pa
et4sv
ett3r
e1tu
etu4ri
et4va
et5vu
e1ty
2etz
e1t^^e4
et^^e4c4
euk4
e5um.
e5up4
4eur
eu4se.
eu5tro
e1v
e4varm
e4vj
ev3r
3exp
ext4r
4e^^e4
f2
3fa
fac4
fac5ke
4fans
4farb
fa3sh
fa4st
fa4t^^f6
4fav
4f3b
f3d
3fe
4fef
fe2l
fes5ta
fe3sto
4fex
2f1f
fff4
ff3l
ff3n
f3fo
ff3r
ffs4
f3f^^e4
ff^^f65re
f3g2
f5h
3fi
fi2br
fib5rig
fi3li
fin5sm
fi3skal
fisk3r
fi2ti
2f3k
1fl
flo4da
4f3m
fma4
1fo
4fof
fol2
folk1
2f5om
fo2na
for4mo
fost3r
4f3p
fra2m
fram5p
f4rer
5freri
fre4s
f4ri.
fri5sp
5frit
fros5ta
fru5str
fr^^e5n5
2f3s
fs2k
f4sl
f4sm
f4sn
f4sp
f4st
f4sv
2ft
f3ta
f4taf
f4tak
f4tap
f4tarm
fte4r
f4tex
f3ti
f4tin
f3to
f4t3r
ft2sa
ft4set
ft2s5i
ft4sj
fts4t
fts5v^^e4
ft5t
ft1v
3fu
furs5te
fu5ru
fu3tu
4fv
5fy
fy4ma
f^^e53t^^f6
1f^^e4
f^^e4s5ti
3f^^f6
f^^f62ra
f^^f62ren
f^^f62ri
f^^f6r3k
f^^f6r3sm
f^^f6r3su
f^^f6rt4
f^^f6r1^^f6
ga5br
3g2ag
4gakt
3g2al
gall3s
ga5l^^e4
ga4no
2garb
4garm
ga2ro
4gart
ga4st
ga4su
5g2ati
gaus4
g4av
g5avsn
4gax
2gb
2gd
g3d4r
ge2a
ge5b4
2gef
2ge4j
g2eli
3gelis
gel5st
gel5y
3gel^^e4
gel5^^e4n
g4em
ge4nap
gen5g
3g2eni
3genj
4genm
genom5
gen4sa
g4ense
1g2ent
4genv
ge5ny
3gen^^e4
ge2o
1g2era
4gerarb
3g2eri
gers5n
5gese
ge4to
get5s
5g2ett
2g1f
2gg
g1ga
g4gap
g1ge
gg5g
gg1l
g4gos
ggs4la
ggs4m
gg3s4t
gg3s4v
g4gu
2gh
gh4te
1g2i
gi1o
gi5sn
gi4ste
gis4tr
gi5stral
gi5st4rat
3giv
gi2^^f6
g2jo
3gjor
g3j^^e4
2g3k2
2gl
g4lans
g1lar
g2las
5glase
glas5k
5glas^^f6
g4lid
4glj
g4l^^f6g
5gl^^f6m
2g1m
2g1n
g4nag
g2no
1g2o
3go.
3gol
gon3s4
4gont
2gord
4gorm
4gort
go3sl
2g1p
g2r4
3graf
5gral
gra2m5
5grans
4gras
5grec
5grett
g3rig
4g5rik
5grip
3gris
g5roi
gro2v
4grum
grus5t
g4r^^e5
5gr^^e5.
gr^^e44n
5gr^^e4ns
2g2s
gs1an
g5satt
g3sel
g4sf
gsi4d
g3sju
g5skaf
gs4ki
gs3kn
gs4kot
g3sky
gs1l
gs1m
g4sme
gs3n
gs4ni
gs4n^^f6
gs1or
gs3pl
gs3po
gs4por
gs5pre
gs3pu
gs3s
gs3tak
gs3tal
g3stark
gs4ten
g3stif
gs3till
gs3tj
g3stol
gs3tra
gst4re
g3st^^e4m
g4sug
gs1v
g4s3ve
gs3vi
gs3v^^e5
gs3yt
gs1^^e4
2g1t
g3tr
1g2u
4gug
guld3
gul4da
4gul^^e4
gu2ma
4gup
gu5ru
gus4k
2gut
g3utb
2g1v
4gw
3gy
gytt3j
1g2^^e5
g^^e5rds5
2g5^^e5ri
g4^^e4l
g2^^e4r
g^^e44s
1g2^^f6
4g^^f6g
g^^f65ro
2g5^^f6rt
1h
ha3bl
ha5ge
ha4li
hal4so
halv3^^e5
ham4st
handels3
hands4l
han5g2a
ha5ra
ha4sc
ha4sp
hasp5l
has3t
hav2
havs3
h5c
4hd
he4at
he4fr
he4l^^e4
hets1
hets3t
hets3v
h3g
h2i
4hir
his2sk
hi4t
hj^^e4l3s
h1k
2hl
h4le
2hm
4hn
h2na
h2nit
ho5nu
hop5plo
hop3s
hos3p
hos5ti
4how
h3p
h5ru
h1s
2ht
hu2s
hust5r
hyg5r
hys4t
hys5ta
hy3ster
h^^e5rd5s4
h^^e4ll2
h^^e4lls1
h^^e4lso3
h^^e44ri
h^^e44s
h^^e44var
h2^^f6
h^^f62g
h^^f65gen
h^^f6g5r
h^^f6rn5s
h^^f64s
h^^f6st5r
i1a
ia3fr
ia3g
ia4lu
ia4sk
ia3tr
i2b3l
i5bril
i3ca
i4ce.
i5cha
ic4kord
ick3u4
i5co
i2d
iden3s
id4ge
i4dom
id1r
id3ro
id2s
ids3v
i4dun
i3d^^e5
i4d^^f6
2i1e
ifes4
i5fn
i1fr
3ifr^^e5n
i1g
4igan
i2geb
ig5ej
ig1l
ig3no
i3i
i4kart
i1ki
i3klo
ik5l^^e4n
ik3n
i1ko
ik3re
i5krob
ik5rof
ik5ros
ik5s2h
ik5skor
i3kul
i3kum
ik5u4t
ik1v
i3ky
i3k^^e5
i3k^^f6
i1la
il4dan
i2lin
il1j^^f6
il5k
il5lak
il4lik
ill3s2
3illu
il5l^^e4r
il2min
i1lo
il2tj
i3lu
ilufts5
i4lup
i5l^^e4
im2b3r
im5sm
im4so
i1mu
i5m^^e5
i3m^^e4
i5m^^f6
i4nau
ind5sk^^e4
ind5sti
1indu
in4ga
in4ge.
ing4es.
ing5is
in5glas
ings5te
i3ni
i4nif
in5j
in5kve
1inneh
5inre
1inri
3inr^^e4
in4sem
in3skr^^e4
in3sl
ins4m
in3sn
1inspe
5inspeln
in5spr
3instink
3instru
in4st^^e5
in5te
1intr
in4tra
int3s
i1nu
i4nun
in3ym
i1n^^e4
i5oc
i1og
i3ok
io4kr
i1ol
io5li
i5om
ion2
i3ono
ions3
i1op
i1or
i1os
i1ot
i1pe
i1pi
ipos4
ip5pi
i3ra
i4res
i1ri
irk5l
i1ro
iro3p
i1ru
i5sce
isel4
is2h
i2sk
is5kep
isk5na
is3kopa
is3ku
is4kun
is3ky
i5slam
is3l^^e4n
is3m
is3n
i2s3p
is4pri
is3sa
is3se
iss5n
is4s3tr
iss3t^^e4
i1stal
i1stans
ist5att
is5ten.
i1stent
is4tes
is3tig
is5ting
is5tor.
is5tore
ist5ro
ist^^e54
is5v
i3sy
i4s^^e5
i1t
it5c
i4tei
i4tex
i4tj
it5ran
i5trin
i3tris
it2t5op
it4t3r
it4tu
i2t5^^e5
4i1u
i1va
i2vak
i1vi
i4vin
iv3r
iv2s
i1v^^e5
ix2t
ix5tu
i1^^f6
1ja
3jakt.
4jarb
jas5p
2jb
2jd
jd3r
jd4sty
j4du
1je
je2a
5jef
je5sta
2j1f
4j3g
4jh
1ji
4jin
4jk
j4kl
j3ko
jk3v
2j1l
2jm
2j1n
j2o
3job
jo4kr
4jolj
jo5l^^f6
jor4din
jord3s4
3jou
4jp
j5pl
2j3r
2j1s
j5sa
j4sk
js4me
js4te
2jt
jts4
2j2u
ju4kos
juk3s
jul3k
4jur
jus5kr
juss4
jus4t
jus5ta
jut4sta
j^^e45lo
j^^e4l4p5r
j^^e4l4sa
j^^e4rn3sk
j^^e4r5s
j^^f6r2s
j^^f6s4t
5j^^e9
1k2a
3ka.
3kad.
3kade.
ka4dr
2kaf
5kaf^^e4
ka3i
ka5ju
2kak
k3akti
4kalf
4kalg
kal4lo
kall3s
3kamp
3kamr
3kan.
4kand.
5kano
2kap
3kapi
ka5pla
kap4pr
kaps5t
5kapten
3kar.
ka3ra
4karb
k5arbet
ka5ri
4kark
3karna
4karp
karp5s
4kart.
4karte
4karv
3kas
ka4sk
kas3ti
3kat.
3kats.
4kau
2kb
4kc
2k3d4
kdom4
1k2e
3ke.
2ked.
2keda
ke3dr
ked4s
ke4er
2kefu
4keld
kels4
4kense
ke5n^^e5
2kep
3kern
ke2s
kes3s
4kex
2k1f
kf^^f62
kf^^f63ri
2k5g4
2kh4
kid3s
4kif
1kig
kik4s
kilt4
5kim^^e5
king3r
4kinne
4kins
2kint
ki4nu
ki4tr
kiv3s
4kj
5kjol
k3j^^e4
2k3k
kl2
1klag
k2lama
kla4mi
3klang.
3klass
2klat
5klav
2kle
k2lej
2klig
k2lim
3klip
k2lis
5klist3r
k5lock.
5klocka
3klos
1klub
4kluk
1kl^^e4d
2k3l^^e4g
2k1m
2k2n
k4nal
3k4nap
5knip
3k4niv
3k4nu
k4ny
k5nyk
k2o
4koc
ko5de
k5odl
kog3n
ko4gr
kog4s3
4kola
ko2lin
4kolj
kol5tr
5kolv.
1kom
3komm
5komp
2k3omr
kom4s
1kon
3konf
3konst
3kont
ko3nu
1kor
3korg
ko3ri
2korr
3korres
5kortera
ko5s4k
ko3sl
3kost
ko4str
4k3ou
2k1p
k2r4
3kraf
5kra3ge
4krang
5krera
k4reten
krid5s2
1krig
krigs3
krings2k
4kriv
3kropp
kropps5
kru5stad
k3ryg
kr^^e5k5s
kr^^e54pa
k5r^^e4dd.
kr^^e4k5l
4kr^^e4l
k3r^^e4t
2ks
ksaks5
k2s5as
ks3ch
k4ser
ks2k4
ks3kl
ks5kra
ks5kv
k3sk^^e4
k3sk^^f6
k5slag.
ks2li
k5sly
k2so
ks3pl
k1s4t
kstavs3
ks5tid
k2su
4k1t
k4tex
kti5ge
k4tinn
k2tins
k2tod
k2tom
k2tr
kt3re
kt3rin
k5trod
kt5rog
kt3rol
kt5r^^e4t
kt2st
kt5t4
k4tug
k2tut
k4t^^e4l
4kug
k5ugn
ku5la
4kuld
3kul^^f6
kum5pl
kungs5
5kunn
ku4pen
ku4ro
3kurs
3kus
kust3a
kv4
3kvali
k5vare
3kvarn
kvar3s
3kvart
k4vato
k2ve
2kvente
1kvinn
5kvire
k4vo
k1v^^e5
3kv^^e4ll
k1v^^e4r
kydds3
ky4lin
3kyrk
k^^e4l4m
5k^^e4mp
5k^^e4nn
3k^^e4ns
3k^^e4rl
4k^^f6g
k^^f6ks5t
5k^^f6p.
k^^f6r4l
k^^f6r4sl
3la.
1lade.
2ladm
4ladr
2laf
3lagd.
la4gin
5lagm
lag3r
2lak
5lakan.
5laki
3laktis
la5lo
3lande.
lan4di
2lappara
2larb
1larn
lar5s
4lart
las3h
4lask
la4st
5laste.
1lat.
la5tr
lat4tis
2lau
2lav
la5vu
2lb4
4l1c
2l2d
lder4s
l3dj
ld3ra
l5dry
lds4an
1le
3le.
le4ge.
le5ig
le2kl
le4kv
lem4s^^f6
2l5enl
3ler.
ler5k
3lern
ler3ste
le5s2l
le5t^^e5
le3um
le4vu
2lex
2l1f
2l1g
l2gj
l3g2l
lgs4
lg5st
2lh
1li
li5ch
3lif
3lig
li4go
lig3s
lik2l
li5kli
lik3s
5limer
2lind
2linga.
ling5o
4lingr
lings5t
2lini
5linj
2lint
li1o
2lip
lis3c
li4sta
li3str^^f6
li4vo
livs1
l2jak
4l1jo
1lju
l5j^^e5
l1j^^e4
l3j^^f6r
2l1k
l3ke
l5kju
l2kl
lk5lag
l5kl^^e4
l2kr
l3k4ra
lk3t
l1la
lld4
ll3dr
lle5b
ll3k
ll1l
l1lo
llok5v
ll3p
ll4san
ll2se
ll3ska
ll2so
ll4sva
ll4tig
ll3tr
l1lu
ll5un
llust3ra
ll5v
l5ly
ll^^e4ggs5
l5l^^f6d
ll^^f6r4
ll5^^f6rt
4l1m
l4mol
lm3st
l1n
lo2af
loc4ku
4lodl
lo4do
lod3st
lo2ge.
2lolj
2lom
4lord
2lorg
lor4s
lo4vo
l4pak
l1pe
l1pi
l5pla
lp5l^^f6
lp4st
4l3r
2l1s
l2sc
l4sjo
l4sj^^e4
l2sk
l4skensv
l3ski
lsk3n
l5skot
l3skr^^e4
l3sky
l3sk^^e5
lsk^^e54p
l3sk^^e4
l3slu
l4sm
ls4mo
ls5nyt
l2sp
l3spe
ls3pl
ls3pol
ls5s
l2st
l3sta
l4stak
ls4te
ls5ter
l3sto
l3sty
l4styg
l3st^^e5
l3st^^e4
l5st^^f6
l2su
l5sur
l2sv
l4svi
ls5vid
l4s^^e5
4l1t
lta2tu
l4tef
l4tif
l4tih
l4tos
lt5rati
l4tret
l4tr^^f6
lt5sk
ltu4
lu5i
luk4to
4lull.
2lun
lung3
2lupp
lu4pu
lus2s5p
5lust.
4lutb
4luts
2lv
l1va
l4varm
lvers4
l1vi
l4vos
lv3ri
lv3sp
l1v^^e4
lv^^e4v4
lycks5t
ly4gat
lyg3r
lyg3s2
3lyste
5lystn
ly4str
2l^^e5.
l^^e5g3s
1l^^e5ng
l^^e5ng3s
l^^e54sk
l^^e5s5te
l^^e54st^^e5
4l^^e4c
l^^e4g5r
1l^^e4nds
5l^^e4ngder
l^^e44san
l^^e44sp
l^^e4tt3s
4l^^f6l
4l^^f6m
3l^^f6n
3l^^f6rer
1l^^f6s
l^^f64v^^e4
3l^^e9
1ma
ma5fr
mag5n
mag5s
ma5ju
mak3r
ma3li
mand4
mang2a
man5g4o
ma5ni
mani1k
5ma3ri
mash5
mas3ko
mask3ro
ma5sk^^f6
mas3ti
mas4v
2mb
mb4sk
2mc
2md
m4dat
m4di
m4do
m3d4r
1me
2meds
me4du
me4kl
me4ko
4meld
melo5
me5lu
men5k
me5nu
me5ny
mer2sko
me4so
mes4t
me3sti
2meta
me5trin
met3ro
meu4
2mex
2m1f
m4fes
m4fn
2m1g4
2mh
1mi
mid3s
mi4lu
2mind
ming4o
4mink
min4kr
4minv
mi3n^^f6
mis2
mi5sf
mi4sp
miss3t
mi4te.
mi4tr
mitt3s
2m1k
2m3l
2m1m2
mme5d
mm3s4
m4mul
2m1n
m2nam
mnas3t
m4nav
mn5dr
mn3g4
mn5st
mn5tu
m2n3^^e5
1mo
m4od
mo4i
2momr
mo3na
mos3k
mo2ta
mo4tin
mo4tu
mot3v
2m1p
m2pak
m4part
m2pl
mp3lad
m5plane
mp3lat
mp3lin
mpos4
mp5p4
mps4k
mp5sp
m4p^^e5
2m1r
4ms
m4sal
m4ske
m3slag
ms3l^^e4
ms2m
mste2
m1sto
m2str
mst3rin
ms5^^e4p
2m1t
4mud
mulls3
mult5r
5mum
4mun3g4
mun4ko
3mur
3musi
mu3sta
mut4sl
2m3v
1myn
mys4te
m^^e5g4
1m^^e5l.
5m^^e5let.
5m^^e5n.
4m^^e5r
m^^e51s
4m^^e4g
m^^e4k3
1m^^e4n
m^^e4ns4
3m^^e4rk
1m^^e4s
m^^e4s5ta
1m^^e4t
m^^f64bl
m^^f64gen.
3m^^f6j
m^^f6r4kl
3m^^f6s
4m^^f6v
1na
3na.
3nad
nads3
2naf
na5gr
2nak
3nako
3nakr
na3kro
n1akt
2nalf
5nalfl
4nalg
nal3s
na2lu
n5amb
5namn
4nand.
4nanv
na4rap
2narb
2nark
4narm
2nart
nast3r
2nb4
2n1c
n2ch
n3cha
n3che
n3chi
ncis4
ncyk3l
2nd
n4dak
n4dav
nd3d4
n5de
nde3s
n4dil
nd5rak
nd5ras
nd3rat
nd3ri
n5dril
n3drop
nd5ros
nd5skal
nd3sn
nds3or
nds5v^^e4
nd5^^e5s
1ne
3ne.
ne4di
5nedl
ne4d3r
ned3s
ne4d^^f6
ne2gr
ne5gres
4nek.
ne5ly
4nenl
ner5sm
nes3s4
ne4sta
ne5s4ti
ne3tre
ne1ut
2nex
2n1f4
nfalls5
nfis3
2ng1
n4gar
n4gen.
n4gend
n4gens
n4genti
n4germ
n4get
n2gi
ng3ig
ngi4s
ng4ly
n2go
ng5om
ng3or
ng3rad
n4gr^^f6
ng4ser
ngs1k
ngs3pa
ngs5tim
ngs3val
n4g^^f6d
2nh
1n2i
4nid
ni5ec
ni4ki
ni5li
3nin
nings1
nings3k
nings5v
ni1o
4nip
nip4pr
ni5steri
nist3ra
ni3t4r
niv5sk
niv5st
2n1j
n4jar
n3jun
nju4s
n3j^^e4
2nk
n4kart
n1ki
n4kis.
n3kny
n1ko
nkrafts5
nk3ri
n1kro
nkrus4
nk5sl
nk3sp
nk4tin
n1ku
n1k^^f6
2n1l
2n1m
2n1n
nn3d
n3ne
nnis4
nn3k
nn3s4t
1no
2nodl
no4kl
2nolj
2nomr
nom3s4
2nord
2norg
no5sa
no5sc
no4tu
2n1p
2n1r
4ns
ns2i
n4sint
n4sis.
n4sise
ns2k
ns3kan
n1ski
ns3kor
nslags5
ns5las
ns5mit
n4soc
n1spi
ns3pl
ns3po
ns3s4
n3stans
n3stap
ns4tel
n3stif
ns3tig
ns4tra
n2strik
nst5up
nst5vil
n3s4ty
n1sva
ns3vi
ns3v^^e4r
2n1t
n4tark
nter5s4
n4tinf
n2t5omb
nt3rad
n3trah
n3trak
n5trala
nt3rali
n5tram
nt3rep
n3trer
nt3ria
nt3rin
nt3ris
n4tropin
n4tror
n4tr^^f6
nts3c
nt4se
nts5kor
nt4str
n4tut
n3tv^^e5
nufts4
4nug
n5ugn
3nui
3num
nums5
2nup
n3upp
2nutb
2n1v
ny5gr
n5z
4n^^e5r
4n^^e4.
4n^^e4c
3n^^e4m
3n^^e4t
4n^^f6g4
3n^^f6j
n^^f62ja
n^^f65kr
4n^^f6l
n^^f6s4
n^^f6s5ke
o1a
o2ard
o2b
5o4bj
o4bli
oby4
oc4k5r
ock3sk
oc3ku
o2d
ode4k
odi4a
1odli
o5dral
o3dro
ods4k
od2st
ods4ti
od5stu
o3d^^e4
o1e
offs5t
o4fl
o3fr
of^^f6rm^^e54
o1g
o4gav
og3gr
o4gj
o5glo
o5gly
ognos4
ogno5st
o4gri
o4gr^^f6
og3se
og4s3t
o4g^^e4
o1i
o4il
o1j
o1k
o4kli
ok3n
ok3sl
ok4su
o2kv
o1la
o5lak
ol5au
olf^^f64
1olj
ol3ka
olk3r
ol4ku
ol4k^^e4
oll4si
oll5sl^^e4
ol3l^^e4
olm4s
oln3s
o1lo
olo5kv
ol4sa
ol4t^^e5
o1lu
o4lug
o4lur
o1ly
ol5^^e5r
o1l^^e4
om4br^^e4
o3men
o4mord
om5pa
om3pl
1omr
4omra
om1sk
om4ste
3oms^^e4t
om4tr
om3tv
on3c
on5gi
on1gr
ongs4l
o4nins
on3j
on1k4
ons3c
onsi3s
ons3m
on5stel
ons4ter
on3tras
on4tre
ont4s
o1ny
on5^^e5
o1n^^e4
o3n^^f6
oo4d
oom5s
o3or
o1pe
o1pi
o5pline
op4pl
opp3le
op4pr
op4pu
o3pri
op4st
o3p^^e5
o5q
4ora
o3rak
oran3g4
o2rap
1ordn
or4d5^^e4
o4reh
1orga
5organi
or4gr
or4g^^e5
o1ri
3orient
4ork
or4m^^f6
or4nu
or4n^^e4
o1ro
or4pl
or5pr
or4spa
ors5tig
or5te
or2tr
ort3re
ort3ro
o1ru
o3ry
o1r^^e4
o1r^^f6
o3s2f^^e4
osk4l
o1skop
o3som
os5pig
os4sk
os4s4t
os3tig
os5tiker
o5still
os4tr
ost5ron
ost5r^^f6
os3tul
ota2lan
4oti.
4otie
4otin
o1to
o5tro
ot5run
ot3sv
ot5ti
ot4tr^^e4
ott2s
o1tu
o5tun
otvin4
o1ty
o5t^^e5
o3t^^e4
oun4
oup4
4our
ou3r^^f6
ou4s
o3ut3t
o1va
ova4n
o1vi
ov3r
ov4si
ov3sl
ovs4me
o1v^^e4
o3we
ox5
oy2
o3^^e5
o3^^e4n
o3^^f6
1pa
4paf
pag4
paki3
pakis4
pa5la
pals5
pa5l^^e4
4pand.
pan4tr
3pap
2parb
4parm
par3s
2pask
pa5ski
pa2st
3patr
pa3u
2pb4
2pc
2p3d4
pek5tri
pekt3ro
4peld
pel3s4i
4pem
5peng
3penn
pent5r
per4bl
3perio
3pers
per4sl
pe5tro
4pex
2p1f
4p3g
2ph
pi4el
1pig
pi1o
3pip
pi5so
pi5sta
pi5sto
p2j
3pj^^e4s
4p3k2
p2l
p4lac
5plan.
p4lane
p3larn
p3lev
3plex
3plic
1plik
4plit
p3lj
1plom
p3lop
2p1m
4p1n
p3ni
1po
5poa
2poc
2pof
po2i
3polit
4polj
poly3
2porg
3pos
pos4ter
4pov
po4v^^e4
2pp
p4part
pp5ask
p4pax
p3pe
p1pi
p4pins
pp3j
pp1l
pp3la
pp3lin
pp5lis
pp5lu
pp3ly
pp3l^^e5n
pp3l^^e5t
pp3l^^e4
pp3l^^f6
pp5oc
pp3of
pp3p4
pp1r
pp3ra
pp3ri
pp3ru
pp3ry
pp3r^^e4
pp3tr
p2pu
p5py
pp3^^e5
p2r2
2pra
5prax
1pres
pres4t
pre3sta
pres5to
p3rig
p3rik
5pril
3princ
pring3
p5riol
3pro
pro3g
p3ror
4pr^^e5
3pr^^e4s
3pr^^f6v
2ps
p2sal
3psalm
p5s2ho
ps4ken
ps2li
p3sna
4pso
p3sod
p1s4t
p4stak
p4st^^e4v
p2s^^f6
2p1t
p3tri
1pu
4pug
pul2l5ov
pul5tr
5pung
3punk
pus3t
2p1v
p^^e53dr
3p^^e4l
p^^e45ro
4p^^f6r
3p^^e9
qu4
3que
1ra
3ra.
raci4t
3rade.
4radr
ra4du
5ra1e
2raff^^e4
ra3fr
ra5is
2rak
ra2lo
r4ande
3rande.
4ran4d3r
rand3s
2ransv
ra3pl
3rar
r4ar.
4rarb
r4are
4rarg
r4ark
4rarm
r4arn
r4ars
4rart
r3arta
ra5r^^f6
r4as
ras3h
ra2st
3raste.
3rativ
ra3tri
2rav
ra5yo
2rb
2r1c
2r2d
r4daf
rda5gr
r3dj
r4dos
rd3ran
rd3rat
r4dul
r3d^^e5
r3d^^e4
r4d^^f6s
1re
3re.
4reaus
re3b
4rec
5reco
re3d4r
re5du
4reft
4regg
3regn.
re1kr
rek5tri
4reld
re3lu
rem5p
3rems
r4en.
2reni
2renk
2renl
re3n^^f6
re3o
3rer.
3rern
3reso
ress5k
re1sti
3ret.
4retet
ret3ro
4rety
re5t^^e5
2revig
4rex
2r1f
rf^^f63ri
2r1g
rg3g2
rgs5top
2rh
rhands5
3rial
4rib
3rifi
2rifr
r3ifr^^e5
3rifu
3rigt
rik2s
3riktn
ri4mo
2rind
rind3s
5ringen.
ring3r
2rinr
2rins
2rint
ri1o
3riot
ri5ple
ri2st^^e4
ri4tut
ri4vis
riv3s
4rj
r4jis
r3jo
r5ju
r5j^^f6
2rk
rk3akt
r4kek
rkes3
r1ki
r3klas
rk2le
r4kl^^f6
rk3n
rk4ne
r1ko
r4kod
rk3tr
r1ku
r4kup
r1k^^e4
r5k^^f6r
2r1l
r5laka
r5lav
rld2
rlds3
rl5sp
2r1m
r4marb
r4mil
rm2s5j
rm5tr
2r1n
rnal4
rn3g4
rn1k
r2nom
rns4k
rns4t
rn3t
ro3b
ro4gro
ro2kr
2rolj
rol4li
rom4a
5roman
5ronau
5rond.
ron4v
ro3pl
ropp2s
ro4ra
2rord
2rorg
2rorie
3rorn
ro4sin
ro4sn
ros3v
ro5te
2r1p
r4pl^^f6
r4p^^f6
4r1r
rra4n
rrd4
rreligi5
rres4
r5rib
rr5k4
r4rob
r4rom
rr1s
rrs2k
r4rur
2rs
r4seld
r4sex
r2sin
r1ski
r4skid
rsk3na
rs5koll
rs4kos
rskotts3
r2sku
r3sk^^f6
rslags4v
r4sle
r4slo
r4s5l^^f6
rs4mo
rs5nat
rs5n^^e4
r1sp
r2spl
r2spo
rs3s4
rs5tak
rs4te
r5stek
rs5tend
r5steni
rs5till
r1sto
r4ston
rst4r
r3str^^f6
r3stu
r1sv
rs4vag
r2sv^^e4
r1sy
2r1t
r2taf
r2takti
rt4an
r4tins
r4tom
r5trit
r3tr^^e4
rt3t
r4tut
rubb5l
ru3br
ru4dan
ruks1
ruks3v
5rullera
3rum.
runn2
runns5
4rupp
rus2h
ru5sha
2rut
5rutig
rut4ra
ru4vi
5ru^^f6
2r1v
rv4sj
rv2s5k^^e4
r3w
rydd5s
ry5o
r^^e5ge5l
4r^^e5l
r^^e5ng3s
r^^e55ra
r^^e53st
r^^e4ck5s
4r^^e4kt
4r^^e4m
r^^e4ng3s
r^^e4ns5t
4r^^e4s
r^^e44san
r^^e4s3s
r^^e45sti
r^^e4v5s
r^^f6d5el
r^^f6d5r
r^^f6d3s
2r^^f6g
r3^^f6i
r^^f6k3s
r^^f6ns4t
4r^^f6p
3r^^f6r
r^^f6r4s
r^^f64st
r^^f6st3r
r1^^f6vr
1sa
3sa.
3sad.
3sade
4sadj
2sa3dr
sad5s
2saf
sa3i
sak5ri
2s1akt
sa5lo
3s2am
sa2ma
samman3
sa2mor
sand3s
4sang
2sanl
s3anl^^e4
san3sla
2sap
3s4ar.
2sarb
2sarm
s5arm.
3sarn
2sart
4sarv
4sass
5sat.
sa4tu
2sau
s3auk
2s1av
4sb
s2c
2sch.
1scha
2schau
4schb
1schen
1scher
1schet
1schi
4schk
4schm
4schp
3schy
3sch^^f6
sci3p
4s3d
1se
se4at.
se2g
2s3egg
3segl
seg3ra
sek5le
sek3r
sek5tr
3sel.
se5ly
sem2
3sen.
s5ers^^e4
3set.
2sexp
2s1f
s4f^^e4r.
sf^^f62
4s3g2
2sh
5s2haw
shi1s
s5h^^f6
1si
sid5s
5sie
si4eri
si4esk
si2ett
3s2ig
3sik
sikts3
5sill.
silver3
silv3r
2s1ind
2s1inf
sinne2s3
3sinni
4sinr
2sin1s
s1inst
5sint.
2sintr
3sio
sis4t
siu4
1s2j
2sjak
s3jakt
4sjn
4sjt
s4ju
5sjuk
4sjur
sj^^e4ls3
3sj^^f6
4sk.
2ska.
3s2kada
s2kado
3skaffn
1skaft
s4kag
s2kal
3skal.
1skap
5skap.
5skapet
4skapi
skaps1
4skar
s4kara
5skarv
4skas
s2kat
s4kav
4ske.
3sked.
s4kene
3skepp
4skh
sk4i
3skif
5skin
4skis.
5skiv
5skjor
3skju
4skl
sk5lap
s3klas
4skn
3s4ko.
1s4kog
4skogsg
1skol
3skola
s4kolo
s4korp
skor1st
1skot
s5kran.
3skrat
sk4ret
3skrev
1skri
3skrif
s3krig
5skrin
3skrip
s5kris
3skriv
s5kron
s4kru
5skrub
3skruv
5skr^^e4c
sk3s
2skt
3skulp
s3kup
2skv
s4kve
1s2ky
s4kyn
2skyrk
1sk^^e5
s4k^^e5l
5sk^^e5p.
4sk^^e5r
5sk^^e4nk
3sk^^e4rv
2sl2
4sla.
s5lad.
s3land
3s2lang
s4lant
s3lar.
4slas
s1lat
s2lev
3slev.
s4lic
slins3
4slis
s2lit
s5lor
slotts3
s2lu
s3luc
s3luf
4slus
s3lust
3slut
slu4to
3sl^^e5.
5s4l^^e5r
s4l^^e4k
s5l^^e4m
s5l^^e4nn
3s4l^^e4p
4s3l^^e4r
s2l^^e4t
3s2l^^f6j
2sm
s2mak
3smak.
s3makt
s2mal
s2met.
s2mid
s2mit
3smitta
s3mj
5smug
5smyg
sm^^e55g
sm^^e53k
sm^^e53s
3sm^^e4d
3sm^^e4l
4sm^^e4s
3sm^^f6r
2s2n4
3snab
3s4nac
s3nam
s5nare
s3nast
s5ner
3snib
3snil
3snit
1snitt
s3niv
3snut
s4n^^e5
5sn^^e5r
5sn^^e4c
s4n^^e4r
3sn^^f6.
sn^^f65g
3sn^^f6r
sn^^f63s
1so
3soc
5sock
2sod
5soi
2solj
sol3s2
2som
5somm
3son
son4st
so5pra
so4pu
3sor.
2sord
s5ord.
2sorg
3sorn
3sot
4sott
s2p2
5spann.
s4park
5sparv
4spas
s3pass
spa5tr
1spe
4sped
3s4pek
3s4pel
4spelsl
2spen
2sper
5spets
3spill
3spir
4spl
s1pla
s3plan
s3plats
spli4
s4plin
5split
s5pl^^e4
4spre
s3pres
4s3pris
3sprit
2spro
s3pry
3spr^^e5
5spr^^e4n
s3ps
1s4p^^e5
3sp^^e5n
3sp^^e5r
5sp^^e4n
3sp^^f6
4s1r
4s1s
s5sad
sse4lin
s5sil
ss2k
ss5kl
ss3kun
ss1l
ss2lag.
ss2l^^e4
ss2l^^f6
ss3na
sss4
ss3unn
s2sv
ss3vi
s2t
2st.
4sta.
5stac
3stadi
s4taf
5stalgis
3stalla
2stalli
5stam.
5stamm
1stant
5stark.
5startad
1state
3statl
1stau
st3c
2s5te.
4stea
5steg.
s4tek.
2stekn
5stekt
s4tell
3stem.
3steme
5stenar
3s4tene
3stense
5stensm
1stera
1stering
s4teriu
3sterne
5stetis
2stia
2stib
3stick
2stid
s4tiken
2stil
3stil.
3stink
3stisc
1stit
2stj
s5tju
3stj^^e4l
3stj^^e4r
2stm
5stoc
1stol
4stolk
4stom
stori4eu
5storis
stor3s
3straff
4strativ
3strato
3strec
3strej
st3ren
1strer
2stria
1strid
5stride
2striel
st4rif
1strikt
st5risk
1stru
3struk
2strumm
s3tryc
5stryk
5str^^e5k
3str^^e5l
3str^^e4c
4str^^e4d
3str^^e4ng
5str^^e4v
3str^^f6m
2st3s4
st3t
4stv
s3tvis
1sty
2styp
1st^^e5
4st^^e5g
5st^^e5l
1st^^e4
3st^^e4l
1st^^f6
1su
su4b
3sug
su3i
3sum
2sun
5sun.
s1under
5sune
s5ung
2sup
5supa
su2pu
5sus
2s1ut
su4to
su4tr
s2v2
5svag.
s3vagn
4s3vak
5svam
4svap
svars3
3svart
4svas
s3vat
4svec
3sven
5svep
4s3ver
s5ves
4s3vil
s4vine
4svis
s5vitt
s5v^^e5d
3sv^^e5ri
3sv^^e4ng
5sv^^e4rm.
s3v^^e4s
s3v^^e4t
4syk
5syl
3syn
syn3k
s3yrk
3sys
sys4t
sys5ter
syt2
sy5th
1s^^e5
5s^^e5g
4s^^e5k
2s^^e5lde
s^^e5ng3
1s^^e4
s4^^e4d
2s5^^e4gg
s4^^e4l
2s^^e4p
5s^^e4s
3s^^e4t
4s^^e4ta
1s^^f6
4s^^f6d
2s^^f6g
s5^^f6ga
s^^f64ko
4s^^f6l
4s^^f6p
s^^f6r2s
2s3^^f6rt
1ta
3ta.
ta1ch
3tade.
4tadi
4tads5
2taff
3taga
5tak.
ta5kre
2taktig
tak4to
4talf
5tallise
tall5s
4talv
3tame
3tami
3tan.
ta4nab
3tande.
2t3anfa
4tanl
t4ap3l
2tappar
3tar.
4tarb
tar4mi
3tarn
tars4
4tart
5tartavl
4tarv
4task
3tast
ta1str
tat2
ta4tan
tats3
2tatt
2tav
4tave
5tavla.
3tavlan
3tavlo
tav2s
3tax
2tb4
2tc
t3cha
t3che
2t3d4
3t2e
te4as
te3b4
5tec
4teg
te2g1r
te3gre
te3i
te4int
4tej
tej2s
te4kl
5teknik
5teknis
4teld
5te5l^^f6
5tema
4temo
te4mu
ten3g4
5tensi
ten3tr
te4n^^e4
te5n^^f6r
5ter.
5teri^^f6
ter3k4
5term
5terna
5ters
ter3t
te4ru
5tes.
5test
tes4te
te5stik
te5stu
5tetik
tets3
4texa
2texp
2t1f4
2t3g4
2th
t4hen
1ti
3tial
5tib
5tici
3tid
5tide
ti4du
4tid^^f6
ti4ed
tifts5
ti2gel
3tigh
ti4go
ti2gr
3tigt
tik3l
3tiks
5tikul
t2il
5tilj
3tillst
3tillv
3till^^e4
5time
2tind
2tinr
2tint
ti4od
3tion
ti2os
3tis
4tisc
5tisk
3tiva
ti4van
5tivite
ti2^^f6
t2j
4tje
4tjob
2tjou
4tj^^e4l
4tj^^e4m
3tj^^e4n
2t3k2
2t3l
2t1m
2t5n4
tne4r
4todl
3tok
4tol.
4tolj
2tomr
4toms
t2op
5torap
t5ord.
5toriett
4torm
torm3s
3torn
tor1st
4tort.
tos4k
t5ost.
t4ov
2t1p
t2r4
2tra
t4raf
3trafi
3t4ral.
t4rala
3t4rale
5tralo
3trals
t4ralt
3trans
tran2s5a
4trar
t3ras.
t3rat.
t4rato
4treg
4tren
4trer.
4trern
t3rets.
2tri
3tribu
5trick
trids3
t5riel
t1ring
t3ring.
2troc
t3rock
t4rog
t5ronik
t3rono
4tropi.
5tross
5trotn
t4rump
t4rup
3trupp
trus5ta
1tryc
5tryck.
5tryggh
4tr^^e5k
5tr^^e4.
3tr^^e4d
tr^^e4ds4
3tr^^e4f
3tr^^e4g
4tr^^e4k
t3r^^e4kn
t4r^^e4n
5tr^^e4ni
5tr^^f6ja
t4r^^f6t
5tr^^e9
2ts
t5s4and
ts5art
t3s4at
t3se
t4seg
ts4en
t4sex
ts2k
t5skall
t3skatt
t1ski
ts3kl
tskotts5
t5slot
ts5l^^e4k
ts3n^^e4
t3sn^^f6
t2so
ts3ord
ts3pl
tss4
t1st
ts4te
ts5ter
ts5tillf
ts3tj
t3stol
t4ston
t2stra
t4stry
t4stur
t5styr
t2su
t3sud
t5sy
2tt
t3tac
t4tau
t4ted
tte5g4
t4tem
tte2n
ttes4
t4tex
t4tins
t4tip
tt3ja
t1to
tt3rad
tt3rand
tt3rat
tt3re
tt3ri
tt4ry
tt4se
tt2si
tt4sta
t3tu
t4tug
tt1v
tt4v^^e5
t3ty
t3t^^e4
t3t^^f6r
4t5ugn
2tund
3tunga
tung3s
5tunn
2tupp
tu5re
2tutb
t3utv
t3ut^^f6
tu4vu
5tu^^f6
2tv
t1va
4tve
t3vig
3tving
t3vit
3tviv
t3v^^e5g
3tv^^e5n
t3v^^e4n
tv^^e4r3s
3tv^^e4tt
ty5da
5tyg.
3tyngd
3typ
ty3pi
5tys
2tz
3t^^e5g
t^^e5s4
4t^^e5t
t^^e4c4ko
4t5^^e4g
4t^^e4m
4t^^e4rm
3t^^e4vl
4t^^f64d
t^^f65de
4t^^f6g
4t^^f6p
t^^f64pi
3t^^f6rer
t^^f6rs3t
t^^f64vas
5t^^e9
u1a
u2b
ub5al
ubb4le
ub3lic
u4bo
u3cha
u5cl
u2d
u4dak
u5de
ud3r
ud4ret
uds4a
u4du
u4dy
u1e
u2es
uf4f^^e4
uf4tan
uf4to
4u1ga
u1ge
ugg3s
ugn4
ugns5
ug3s4
u5ie
u1in
u3is
u3itet
u3j
u2keb
u5ki
u4kl
uk5la
uk3n
u1ko
ukos4
uk2s
uks5ko
uk3tris
ukt5s
uk4t^^e4
u3ku
uk3v
u1la
ul4di
ulds2m
ul4du
ul4d^^f6
ull3ste
ull3^^e4n
u1lo
uls5ti
ul2tr
u3lu
u1l^^e4
u1l^^f6
um4f^^e4
um4so
ums4t
u1mu
u3m^^f6r
5underl
1unders^^f6
1underv
un4dom
und3r
un4d^^e5
un5g2ef
un3gersk
ung5it
ung3r
ungs4p
3unif
unk3l
unk3n
un4kr
un1sk
un4tr
un5trati
u5nu
u1o
u1pe
u4pern
u1pi
u2pl
u3plet
up3lik
3uppfa
1uppg
up4pin
1uppla
5uppl^^e4
up4p3r
upp3s
upp5sp
up5ut
ur5ak
ur5arv
u3re
u1ri
u1ro
u4rob
u4rom
urs5tin
ur4st^^e4
u5ry
u2sak
us5anl
u3scha
u3se
usen3
u2s1k
us3ka
us4kla
us4kr
u5sky
us4k^^e5
us5l^^e4
us3n
u2sp
us3pen
us5tat
us3tig
u3stik
us5tin
ust5ro
u4st^^e5
u4st^^e4
us3v
u4s^^e5
u4s^^e4
u2s^^f6
u4tak
1utb
u4tef
ute3s
utik2
u5til
uti3^^f6
ut3j
3utj^^e4m
utlands3
u1to
u3top
uto5s
ut3r
ut4rer
ut4ro
ut5rop
1utru
2utsid
ut3sl
3utsl^^e4
2utt
utt4j
ut1v
3utvec
u5ty
ut3^^f6v
u5u
2u1v
u2vak
u4vj
u4v^^e4
u5^^e5
u3^^f6
va5dro
1vagn
2v1akti
val3k
val4li
val4st
5valv
5vama
4vand.
4vanp
van4st
van5tr
5vap
2varb
va4res
va4ri.
4vark
var2s
vart5r
va1ru
vas5ti
5vattn
4vau
4vav
5vavi
2vb4
2v1c
2v3d4
1ve
5vec
ve2k
ve3ke
4veld
vensk3^^e4
5ventera
ve3ny
ve5n^^f6
4vep
ver5g
3verk
ves4
ve2s5p
ve1st
3veta
3vete
vet5sa
vett5s
2v1f
2v1g
2vh
v4i
vi4c
vid3s
vild3s
vil4t
3vind.
ving3s4
3vinkl
vi2no
5vinst.
5vinste
vi5ny
3vis.
vi5sa
vis5h
vis5ko
vi4st
vis3ta
vi2tr
vi4var
4vjo
2v3k2
2v1l
2v1m
vm^^f6rk4
2v1n4
1vo
4vok.
2vom
4vord
2vorg
vos4
2v1p
2v2r
5vrak
3vrera
v3ru
2vs
v4sc
v1s2k
v2skri
vs4mi
v3sni
v2so
v1st
vs4te
vs5tr^^e5
v5styc
vs3v^^e5
v2s^^f6
2v1t
vu4d1
v1und
4v5up
4vut
2v1v
3vy
5v^^e5ld
v^^e5ngs3
3v^^e5rd
4v^^e5ri
v^^e53ru
3v^^e4g
v^^e4gg5s
v^^e44l
v^^e4ll4s3
3v^^e4nl
3v^^e4rde
v^^e44ril
4v^^e4rj
5v^^e4rk
3v^^e4rld
2v^^e4t
3v^^e4x
4v^^f6g
4v^^f6p
3v^^f6r
1wa
we2
w2h
whi2
wi2e
w4na
x1
xan5d4
xem3pla
xis4
xk2
xli4
xs4
xti2
x4t^^e5
2y
y1a
y4bris
yb4s
y2d
y4da
y5dan
y4do
yd3r
yds4
y4du
y4d^^f6
y1e
y1ga
y1ge
ygg3r
yg4g^^e5
ygs4p
y1i
y1ki
y5klist
yk5lon
yk3n
y1ko
y1la
yl4gj
y3li
yl5k
yl5l^^e4
y1lo
yl4tr
ym2fl
ym4for
y3m^^e5
yng3r
ynk5l
yn4sa
yns4t
y3or
y5ou
y1pe
y5po
yp3ri
yre4s
y1ri
yr4ku
yrk5v
y1ro
yrs4k
yr5st
yr5tu
y1r^^e53
y5scho
ys2st
ys3ta
ys3ti
ys4tik.
yst3ra
y2tak
y4te.
y4tea
y1to
ytt3r
yt5v
y3va
y3vi
y3v^^e4
y5w
y5^^e5
1za
1ze
ze4ro
1zi
1zo
zo4nal
4zp
z5s
3zu
z4zin
^^e51a
^^e53dj
^^e5ds4l
^^e51e
^^e51f
^^e51ga
^^e51ge
^^e5ge2l
^^e5g3l
^^e5g3s4k
^^e5g3st
^^e5g^^e54
^^e53i
^^e51ki
5^^e5klag
^^e5k4str^^e4
^^e51la
1^^e5lder
^^e52lin
^^e5l3k
^^e5ll4sp
^^e5l2s5e
^^e5l3st
^^e51l^^e4
^^e51m
^^e5man4s
^^e5nd4r
^^e5n4du
^^e5ns4t
^^e5ns4v
^^e53o
^^e51p
^^e52pl
^^e55pla
^^e54p^^f6
^^e5r4do
^^e5rd4ra
^^e5rd2s
^^e5rd4s3t
^^e54rel
^^e51ri
^^e55ror
5^^e5rsav
^^e5r5s2li
^^e5r2sv
^^e5r5^^f6
^^e5s4ke
^^e5s3n
^^e5ss4
^^e5s4skr
^^e5s4t
^^e5te2
^^e5t3ri
^^e53tr^^e5
^^e5t2sj
^^e5tt5s
^^e51v
^^e41a
^^e42b
2^^e4c
^^e4ck5v
^^e42d
^^e4dd3s
^^e4d4du
^^e4de4s
^^e4d3r
^^e4d5se
^^e4d3st
^^e43e
^^e41ga
^^e41ge
^^e4g4go
^^e4g1l
^^e4g3r
^^e4g4re
^^e4g3se
^^e43i
^^e45jo
4^^e4k
^^e41ki
^^e4k3n
^^e4k3r
^^e41la
^^e4l4pap
^^e4l4seg
^^e4ls5kog
^^e4l4slu
^^e4l2t3r
^^e4l2tu
^^e4l4vin
^^e4mp3l
4^^e4ndligh
^^e4nd3r
^^e4nd1st
^^e4ng5r
^^e4nni3s
^^e4nn3s
^^e44no
^^e4ns1l
^^e4n4st
^^e4ns5te
^^e4n4sv
^^e4n2t3r
^^e43pe
^^e4pp3l
^^e44pr
^^e4p4st
^^e44rap
^^e4r2bre
^^e4rg5l
^^e4r4gr
^^e41ri
^^e4rib4
^^e4r4k^^e4
^^e4r4nis
^^e4rn3st
^^e4r2n^^e5
^^e4r4n^^f6
^^e4r5ob
^^e45rol
^^e43rop
^^e45ror
^^e45ros
^^e4r2si
^^e4r4sko
^^e4r2so
^^e4r4sp
^^e4r2sv
^^e4r4tand
^^e4r2tr
^^e4rt3s
4^^e4s
^^e4s3pa
^^e4s5pi
^^e4s4sk
^^e4s4sp
^^e4s3ta
^^e4st3r
^^e44st^^e4
^^e44s^^e5
2^^e4t
^^e43to
^^e45tre
^^e4t4s3k
^^e4t5te
^^e4t4top
^^e4tt3r
^^e4t4tu
^^e4t4tv
^^e41va
^^e42vak
^^e43vi
^^e45vu
^^f61a
^^f62d
^^f64dak
^^f64dal
^^f64darv
^^f6de4s5
^^f64dis
^^f6d3ra
^^f6d2s
^^f6d3se
^^f64du
^^f64d^^f6
^^f61e
^^f61ga
^^f6g5ak
^^f65gar
1^^f6gd
^^f61ge
^^f65ger
^^f6gg4
^^f6g1l
^^f6g2n
^^f6gn3e
1^^f6go
^^f6g3si
^^f6g3sk
^^f61i
^^f63jo
^^f6j4sv
^^f64karm
^^f61ki
^^f6k3n
^^f6k2s
^^f6k3sl
^^f61la
^^f6l4kv
^^f6l4k^^f6
^^f6l2p
^^f65l^^e4
^^f6man4
^^f6m2kl
^^f64nal
^^f62nom
^^f6ns3ke
^^f6n4so
^^f6nst3r
^^f63pe
^^f64pel
^^f63pi
^^f6p5li
^^f65plo
1^^f6ppn
^^f64pr
^^f63rande
^^f63ras
^^f64rask
^^f6rb4
^^f6r3d4r
^^f6r1eni
^^f63res
^^f64restr
^^f63ret
^^f6r5evig
^^f6r3g
^^f61ri
^^f65rig
^^f63ring
^^f6r3int
^^f6r5ir
^^f6r5iv
^^f6r4kal
^^f6r1k2l
^^f6r5kli
^^f6r4nis
^^f6r3ol
^^f6r1or
^^f6r2p5la
^^f6r1s2k
^^f6r3sl
^^f6r4sl^^e4
^^f6r5te
^^f6rt5s
^^f6r1u
^^f6r3vr
^^f6r3y
^^f6r1^^e4
^^f6r^^f64d
^^f62sak
^^f6s3n
^^f6s4sj
^^f6s2sk
^^f6s4sp
^^f6s3ta
^^f6st3v
^^f62tak
^^f6ts5ko
^^f6t4st
^^f61v
^^f6ve4
^^f6ver1
5^^f6vere
^^f62vj
^^f6v3ra
^^f6v3ri
^^f6v4sk
^^e93e
}
}

% s-ts-mode
